magic
tech scmos
timestamp 1594036216
<< nwell >>
rect -17 -10 29 8
<< ptransistor >>
rect -5 -4 -3 2
rect 15 -4 17 2
<< pdiffusion >>
rect -11 1 -5 2
rect -11 -3 -10 1
rect -6 -3 -5 1
rect -11 -4 -5 -3
rect -3 1 3 2
rect -3 -3 -2 1
rect 2 -3 3 1
rect -3 -4 3 -3
rect 9 1 15 2
rect 9 -3 10 1
rect 14 -3 15 1
rect 9 -4 15 -3
rect 17 1 23 2
rect 17 -3 18 1
rect 22 -3 23 1
rect 17 -4 23 -3
<< pdcontact >>
rect -10 -3 -6 1
rect -2 -3 2 1
rect 10 -3 14 1
rect 18 -3 22 1
<< psubstratepcontact >>
rect 0 -27 4 -23
rect 13 -27 17 -23
<< nsubstratencontact >>
rect -14 10 -10 14
rect -4 10 0 14
rect 6 10 10 14
rect 16 10 20 14
<< polysilicon >>
rect -5 2 -3 4
rect 15 2 17 4
rect -5 -12 -3 -4
rect 15 -12 17 -4
rect -5 -14 17 -12
<< metal1 >>
rect -15 10 -14 14
rect -10 10 -4 14
rect 0 10 6 14
rect 10 10 16 14
rect 20 10 24 14
rect -10 1 -6 10
rect 10 1 14 10
rect -2 -16 2 -3
rect 18 -16 22 -3
rect -2 -20 22 -16
rect 7 -23 11 -20
rect -6 -27 0 -23
rect 4 -27 13 -23
rect 17 -27 24 -23
<< labels >>
rlabel polysilicon -5 -14 -3 -11 1 BL
rlabel polysilicon 15 -14 17 -9 1 BLbar
<< end >>
